module InstructionModule
#(

);
